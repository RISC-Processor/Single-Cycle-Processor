moduel ALU (
    input wire [31:0] srcA,
    input wire [31:0] srcB,
    input wire [2:0] ALUControl,
    output wire [31:0] ALUResult
);

assign ALUResult = (ALUOp == 3'b010) ? srcA + srcB ;

endmodule